/*
 * Copyright (c) 2020 The VxEngine Project. All rights reserved.
 *
 * Redistribution and use in source and binary forms, with or without
 * modification, are permitted provided that the following conditions
 * are met:
 * 1. Redistributions of source code must retain the above copyright
 *    notice, this list of conditions and the following disclaimer.
 * 2. Redistributions in binary form must reproduce the above copyright
 *    notice, this list of conditions and the following disclaimer in the
 *    documentation and/or other materials provided with the distribution.
 *
 * THIS SOFTWARE IS PROVIDED BY THE AUTHOR AND CONTRIBUTORS ``AS IS'' AND
 * ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
 * IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
 * ARE DISCLAIMED.  IN NO EVENT SHALL THE AUTHOR OR CONTRIBUTORS BE LIABLE
 * FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
 * DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
 * OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
 * HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT
 * LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY
 * OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF
 * SUCH DAMAGE.
 */

/*
 * Floating point exponent alignment module
 */

module flp_align(
	i_sg1,
	i_ex1,
	i_sg2,
	i_ex2,
	o_sg1,
	o_sg2,
	o_ex
);
parameter EWIDTH = 8;		/* Exponent width */
parameter SWIDTH = 23;		/* Significand width */
parameter RSWIDTH = 2;		/* Reserved width for rounding */
localparam OUTWIDTH = 1 + SWIDTH + RSWIDTH;
/* Inputs */
input wire [SWIDTH:0]		i_sg1;	/* Significand 1 */
input wire [EWIDTH-1:0]		i_ex1;	/* Exponent 1 */
input wire [SWIDTH:0]		i_sg2;	/* Significand 2 */
input wire [EWIDTH-1:0]		i_ex2;	/* Exponent 2 */
/* Outputs */
output reg [OUTWIDTH-1:0]	o_sg1;	/* Aligned significand 1 */
output reg [OUTWIDTH-1:0]	o_sg2;	/* Aligned significand 2 */
output wire [EWIDTH-1:0]	o_ex;		/* Common exponent */


wire [EWIDTH:0]		exd;	/* Exponent delta */
wire			exneg;	/* Exponent delta is negative */
wire [EWIDTH-1:0]	shamt;	/* Significand shift amount */
wire [SWIDTH:0]		shsg;	/* Significand which need to be shifted */
wire [OUTWIDTH-1:0]	sg[0:SWIDTH];	/* Shifted significands */

assign exd = { 1'b0, i_ex1 } - { 1'b0, i_ex2 };
assign exneg = exd[EWIDTH];
assign shamt = exneg ? -exd[EWIDTH-1:0] : exd[EWIDTH-1:0];
assign shsg = exneg ? i_sg1 : i_sg2;


genvar g;

/* Generate right shifts */
generate
for(g = SWIDTH; g >= RSWIDTH; g = g-1)
begin: shr
	flp_shrjam #(
		.INWIDTH(OUTWIDTH),
		.OUTWIDTH(OUTWIDTH),
		.SHAMT(g-RSWIDTH)
	) shift_r (
		.in({ {RSWIDTH{1'b0}}, shsg }),
		.out(sg[g])
	);
end
endgenerate

/* Generate left shifts */
generate
for(g = RSWIDTH-1; g >= 0; g = g-1)
begin: shl
	flp_shlpad #(
		.INWIDTH(OUTWIDTH),
		.OUTWIDTH(OUTWIDTH),
		.SHAMT(RSWIDTH-g)
	) shift_l (
		.in({ {RSWIDTH{1'b0}}, shsg }),
		.out(sg[g])
	);
end
endgenerate


assign o_ex = exneg ? i_ex2 : i_ex1;

`define IDX_WIDTH(x)		\
	(x <= 2) ? 1 :		\
	(x <= 4) ? 2 :		\
	(x <= 8) ? 3 :		\
	(x <= 16) ? 4 :		\
	(x <= 32) ? 5 :		\
	(x <= 64) ? 6 :		\
	(x <= 128) ? 7 :	\
	(x <= 256) ? 8 :	\
	-1
localparam IW = `IDX_WIDTH(SWIDTH+1);
`undef IDX_WIDTH

/* Multiplexing logic depending on shift amount */
always @(*)
begin
	o_sg1 = {OUTWIDTH{1'b0}};
	o_sg2 = {OUTWIDTH{1'b0}};

	if(shamt <= SWIDTH)
	begin
		o_sg1 = exneg ? sg[shamt[IW-1:0]] : { i_sg1, {RSWIDTH{1'b0}} };
		o_sg2 = !exneg ? sg[shamt[IW-1:0]] : { i_sg2, {RSWIDTH{1'b0}} };
	end
	else
	begin
		o_sg1 = exneg ? {OUTWIDTH{1'b0}} : { i_sg1, {RSWIDTH{1'b0}} };
		o_sg2 = !exneg ? {OUTWIDTH{1'b0}} : { i_sg2, {RSWIDTH{1'b0}} };
	end
end


endmodule /* flp_align */
