/*
 * Copyright (c) 2020-2023 The VxEngine Project. All rights reserved.
 *
 * Redistribution and use in source and binary forms, with or without
 * modification, are permitted provided that the following conditions
 * are met:
 * 1. Redistributions of source code must retain the above copyright
 *    notice, this list of conditions and the following disclaimer.
 * 2. Redistributions in binary form must reproduce the above copyright
 *    notice, this list of conditions and the following disclaimer in the
 *    documentation and/or other materials provided with the distribution.
 *
 * THIS SOFTWARE IS PROVIDED BY THE AUTHOR AND CONTRIBUTORS ``AS IS'' AND
 * ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
 * IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
 * ARE DISCLAIMED.  IN NO EVENT SHALL THE AUTHOR OR CONTRIBUTORS BE LIABLE
 * FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
 * DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
 * OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
 * HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT
 * LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY
 * OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF
 * SUCH DAMAGE.
 */

/*
 * Parameterized register with reset signal
 */


/* Register */
module vxe_reg_rst #(
	parameter DATA_WIDTH = 32,	/* Register data width */
	parameter RST_VALUE = 0		/* Reset value */
)
(
	clk,
	nrst,
	/* Write control */
	wr_en,
	/* Data in/out */
	data_in,
	data_out
);
localparam [DATA_WIDTH-1:0]	RV = RST_VALUE;
/**/
input wire			clk;
input wire			nrst;
/* Write control */
input wire			wr_en;
/* Data in/out */
input wire [DATA_WIDTH-1:0]	data_in;
output wire [DATA_WIDTH-1:0]	data_out;


reg [DATA_WIDTH-1:0] q;

always @(posedge clk or negedge nrst)
begin
	if(!nrst)
		q <= RV;
	else if(wr_en)
		q <= data_in;
end


assign data_out = q;

endmodule /* vxe_reg_rst */
